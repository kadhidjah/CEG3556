--------------------------------------------------------------------------------
-- Title         : 3-bit Shift Register
-- Project       : VHDL Synthesis Overview
-------------------------------------------------------------------------------
-- File          : threeBitShiftRegister.vhd
-- Author        : Rami Abielmona  <rabielmo@site.uottawa.ca>
-- Created       : 2003/05/17
-- Last modified : 2007/09/25
-------------------------------------------------------------------------------
-- Description : This file creates a 3-bit shift register as defined in the VHDL 
--		 Synthesis lecture. The architecture is done at the RTL 
--		 abstraction level and the implementation is done in structural
--		 VHDL.
-------------------------------------------------------------------------------
-- Modification history :
-- 2003.05.17 	R. Abielmona		Creation
-- 2004.09.22 	R. Abielmona		Ported for CEG 3550
-- 2007.09.25 	R. Abielmona		Modified copyright notice
-------------------------------------------------------------------------------
-- This file is copyright material of Rami Abielmona, Ph.D., P.Eng., Chief Research
-- Scientist at Larus Technologies.  Permission to make digital or hard copies of part
-- or all of this work for personal or classroom use is granted without fee
-- provided that copies are not made or distributed for profit or commercial
-- advantage and that copies bear this notice and the full citation of this work.
-- Prior permission is required to copy, republish, redistribute or post this work.
-- This notice is adapted from the ACM copyright notice.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY threeBitShiftRegister IS
	PORT(
		i_resetBar, i_load	: IN	STD_LOGIC;
		i_clock			: IN	STD_LOGIC;
		i_Value			: IN	STD_LOGIC;
		o_Value			: OUT	STD_LOGIC);
END threeBitShiftRegister;

ARCHITECTURE rtl OF threeBitShiftRegister IS
	SIGNAL int_Value, int_notValue : STD_LOGIC_VECTOR(22 downto 0);

	COMPONENT enARdFF_2
		PORT(
			i_resetBar	: IN	STD_LOGIC;
			i_d		: IN	STD_LOGIC;
			i_enable	: IN	STD_LOGIC;
			i_clock		: IN	STD_LOGIC;
			o_q, o_qBar	: OUT	STD_LOGIC);
	END COMPONENT;

BEGIN

msb: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => i_Value, 
			  i_enable => i_load,
			  i_clock => i_clock,
			  o_q => int_Value(22),
	          o_qBar => int_notValue(22));

ssb: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(22),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(21),
	          o_qBar => int_notValue(21));
ssb1: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(21),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(20),
	          o_qBar => int_notValue(20));
ssb2: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(20),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(19),
	          o_qBar => int_notValue(19));
ssb3: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(19),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(18),
	          o_qBar => int_notValue(18));
ssb4: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(18),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(17),
	          o_qBar => int_notValue(17));
				 
ssb5: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(17),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(16),
	          o_qBar => int_notValue(16));
ssb6: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(16),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(15),
	          o_qBar => int_notValue(15));
ssb7: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(15),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(14),
	          o_qBar => int_notValue(14));
ssb8: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(14),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(13),
	          o_qBar => int_notValue(13));
ssb9: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(13),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(12),
	          o_qBar => int_notValue(12));
ssb10: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(12),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(11),
	          o_qBar => int_notValue(11));
ssb11: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(10),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(),
	          o_qBar => int_notValue(9));
ssb12: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(9),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(8),
	          o_qBar => int_notValue(8));
ssb13: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(8),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(7),
	          o_qBar => int_notValue(7));
ssb14: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(7),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(6),
	          o_qBar => int_notValue(6));
ssb15: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(6),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(5),
	          o_qBar => int_notValue(5));
ssb16: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(5),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(4),
	          o_qBar => int_notValue(4));
ssb17: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(4),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(3),
	          o_qBar => int_notValue(3));
ssb18: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(3),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(2),
	          o_qBar => int_notValue(2));
ssb19: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(2),
			  i_enable => i_load, 
			  i_clock => i_clock,
			  o_q => int_Value(1),
	          o_qBar => int_notValue(1));
lsb: enARdFF_2
	PORT MAP (i_resetBar => i_resetBar,
			  i_d => int_Value(1), 
			  i_enable => i_load,
			  i_clock => i_clock,
			  o_q => int_Value(0),
	          o_qBar => int_notValue(0));

	-- Output Driver
	o_Value		<= int_Value(0);

END rtl;
